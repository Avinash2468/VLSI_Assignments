`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:56:09 09/26/2019
// Design Name:   CRA
// Module Name:   /home/avinash/Desktop/vlsi_lab3/FA/CRA_test.v
// Project Name:  FA
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: CRA
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module CRA_test;

	// Inputs
	reg [3:0] x;
	reg [3:0] y;
	reg c_in;

	// Outputs
	wire c_out;
	wire [3:0] sum;

	// Instantiate the Unit Under Test (UUT)
	CRA uut (
		.c_out(c_out), 
		.sum(sum), 
		.x(x), 
		.y(y), 
		.c_in(c_in)
	);

	initial begin
		// Initialize Inputs
		x = 4'b0000;
		y = 4'b0000;
		c_in = 0;
		// Wait 100 ns for global reset to finish
		#3.5;
      repeat(15)
		begin
		y = 4'b0000;
		repeat(15)
		begin
		#3.5;
		y = y + 4'b0001;
		end
		#3.5;
		x = x+4'b0001;
		end
		// Add stimulus here

	end
      
endmodule

